module PPUAttributeAddress(
    /* verilator lint_off UNUSED */
    input i_clk,
    input i_reset_n
    /* verilator lint_on UNUSED */
);

// https://wiki.nesdev.com/w/index.php/PPU_scrolling#Tile_and_attribute_fetching

endmodule
